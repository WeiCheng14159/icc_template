module BONDPADCNU ();
endmodule
module BONDPADCGU ();
endmodule
