.SUBCKT BONDPADCNU
.ENDS

.SUBCKT BONDPADCGU
.ENDS
